module thirty_two_bit_alu(a, b, Cin, less, op, R, Cout, V);
input [31:0] a;
input [31:0] b;
input [2:0] op;
input Cin, less;
output [31:0] R;
output Cout, V;
wire C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15, C16, C17, C18, C19, C20, C21, C22, C23, C24, C25, C26, C27, C28, C29, C30, C31, slt;
one_bit_alu one_0(a[0], b[0], Cin, slt, op, R[0], C1);
one_bit_alu two_0(a[1], b[1], C1, 1'b0, op, R[1], C2);
one_bit_alu three_0(a[2], b[2], C2, 1'b0, op, R[2], C3);
one_bit_alu four_0(a[3], b[3], C3, 1'b0, op, R[3], C4);
one_bit_alu five_0(a[4], b[4], C4, 1'b0, op, R[4], C5);
one_bit_alu six_0(a[5], b[5], C5, 1'b0, op, R[5], C6);
one_bit_alu seven_0(a[6], b[6], C6, 1'b0, op, R[6], C7);
one_bit_alu eight_0(a[7], b[7], C7, 1'b0, op, R[7], C8);
one_bit_alu one_1(a[8], b[8], C8, 1'b0, op, R[8], C9);
one_bit_alu two_1(a[9], b[9], C9, 1'b0, op, R[9], C10);
one_bit_alu three_1(a[10], b[10], C10, 1'b0, op, R[10], C11);
one_bit_alu four_1(a[11], b[11], C11, 1'b0, op, R[11], C12);
one_bit_alu five_1(a[12], b[12], C12, 1'b0, op, R[12], C13);
one_bit_alu six_1(a[13], b[13], C13, 1'b0, op, R[13], C14);
one_bit_alu seven_1(a[14], b[14], C14, 1'b0, op, R[14], C15);
one_bit_alu eight_1(a[15], b[15], C15, 1'b0, op, R[15], C16);
one_bit_alu one_2(a[16], b[16], C16, 1'b0, op, R[16], C17);
one_bit_alu two_2(a[17], b[17], C17, 1'b0, op, R[17], C18);
one_bit_alu three_2(a[18], b[18], C18, 1'b0, op, R[18], C19);
one_bit_alu four_2(a[19], b[19], C19, 1'b0, op, R[19], C20);
one_bit_alu five_2(a[20], b[20], C20, 1'b0, op, R[20], C21);
one_bit_alu six_2(a[21], b[21], C21, 1'b0, op, R[21], C22);
one_bit_alu seven_2(a[22], b[22], C22, 1'b0, op, R[22], C23);
one_bit_alu eight_2(a[23], b[23], C23, 1'b0, op, R[23], C24);
one_bit_alu one_3(a[24], b[24], C24, 1'b0, op, R[24], C25);
one_bit_alu two_3(a[25], b[25], C25, 1'b0, op, R[25], C26);
one_bit_alu three_3(a[26], b[26], C26, 1'b0, op, R[26], C27);
one_bit_alu four_3(a[27], b[27], C27, 1'b0, op, R[27], C28);
one_bit_alu five_3(a[28], b[28], C28, 1'b0, op, R[28], C29);
one_bit_alu six_3(a[29], b[29], C29, 1'b0, op, R[29], C30);
one_bit_alu seven_3(a[30], b[30], C30, 1'b0, op, R[30], C31);
one_bit_alu_msb eight_3(a[31], b[31], C31, 1'b0, op, R[31], Cout, V, slt);
endmodule