module extendUpper (upper, result);
input [15:0] upper;
output [31:0] result;
and(result[0], 1'b0, 1'b1);
and(result[1], 1'b0, 1'b1);
and(result[2], 1'b0, 1'b1);
and(result[3], 1'b0, 1'b1);
and(result[4], 1'b0, 1'b1);
and(result[5], 1'b0, 1'b1);
and(result[6], 1'b0, 1'b1);
and(result[7], 1'b0, 1'b1);
and(result[8], 1'b0, 1'b1);
and(result[9], 1'b0, 1'b1);
and(result[10], 1'b0, 1'b1);
and(result[11], 1'b0, 1'b1);
and(result[12], 1'b0, 1'b1);
and(result[13], 1'b0, 1'b1);
and(result[14], 1'b0, 1'b1);
and(result[15], 1'b0, 1'b1);
and(result[16], upper[0], 1'b1);
and(result[17], upper[1], 1'b1);
and(result[18], upper[2], 1'b1);
and(result[19], upper[3], 1'b1);
and(result[20], upper[4], 1'b1);
and(result[21], upper[5], 1'b1);
and(result[22], upper[6], 1'b1);
and(result[23], upper[7], 1'b1);
and(result[24], upper[8], 1'b1);
and(result[25], upper[9], 1'b1);
and(result[26], upper[10], 1'b1);
and(result[27], upper[11], 1'b1);
and(result[28], upper[12], 1'b1);
and(result[29], upper[13], 1'b1);
and(result[30], upper[14], 1'b1);
and(result[31], upper[15], 1'b1);
endmodule