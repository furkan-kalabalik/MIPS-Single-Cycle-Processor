module mips32(result, clk);
input clk;
wire [31:0] instruction;
output [31:0] result;
wire RegWrite, AluSrc, MemtoReg, MemRead, MemWrite, LuiCtrl, LoadCtrl, StoreCtrl;
wire [1:0] ALUop;
wire [2:0] ALUctr;
wire [31:0] read_data_1;
wire [31:0] read_data_2;
wire [31:0] singExtendResult;
wire [31:0] registerOutputMux;
wire [31:0] ALUResult;
wire Cout, V;
wire [31:0] memReadResult;
wire [31:0] extendUpperResult;
wire [31:0] selectedResult;
wire [31:0] lbRes;
wire [31:0] lhRes;
wire [31:0] lbuRes;
wire [31:0] lhuRes;
wire [31:0] load4x1Result;
wire [31:0] loadResult;
wire [31:0] sbRes;
wire [31:0] shRes;
wire [31:0] store2x1Result;
wire [31:0] storeResult;
program_counter pc(instruction,clk);
ControlUnit test2(instruction[31:26], RegWrite, AluSrc, MemtoReg, MemRead, MemWrite, ALUop, LuiCtrl, LoadCtrl, StoreCtrl);
ALUCtrl aluCont(instruction[5:0], ALUop, ALUctr);	
extendUpper extend(instruction[15:0], extendUpperResult);
muxTwotoOne32Bit selectResult(loadResult, extendUpperResult, LuiCtrl, selectedResult);
mips_registers registers(read_data_1, read_data_2, selectedResult, instruction[25:21], instruction[20:16], instruction[20:16], RegWrite, clk );
signExtend16Bit ext(instruction[15:0], singExtendResult);
muxTwotoOne32Bit registerOut(read_data_2, singExtendResult, AluSrc, registerOutputMux);
thirty_two_bit_alu ALU(read_data_1, registerOutputMux, ALUctr[2], 1'b0, ALUctr, ALUResult, Cout, V);
extend8BitSigned sbextend(read_data_2, sbRes);
extend16BitSigned shextend(read_data_2, shRes);
muxTwotoOne32Bit selectSW(sbRes, shRes, instruction[26], store2x1Result);
muxTwotoOne32Bit selectStored(store2x1Result, read_data_2, StoreCtrl, storeResult);
mips_memory mem( memReadResult, storeResult, ALUResult, MemWrite, MemRead, clk);
muxTwotoOne32Bit memOut(ALUResult, memReadResult, MemtoReg, result);
extend8BitSigned lbextend(result, lbRes);
extend8BitUnsigned lbuextend(result, lbuRes);
extend16BitSigned lhextend(result, lhRes);
extend16BitUnsigned lhuextend(result, lhuRes);
mux_4x1_32Bit loadHalfOrLoadByte(instruction[26], instruction[28], lbRes, lhRes, lbuRes, lhuRes, load4x1Result);
muxTwotoOne32Bit loadedVal(load4x1Result, result, LoadCtrl, loadResult);
endmodule