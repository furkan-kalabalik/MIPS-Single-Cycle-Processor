module mux_4x1_32Bit(S0,S1, I0, I1, I2, I3, R);
input [31:0] I0;
input [31:0] I1;
input [31:0] I2;
input [31:0] I3;
input S0, S1;
output [31:0] R;

mux_4x1 one(S0,S1, I0[0], I1[0], I2[0], I3[0], R[0]);
mux_4x1 two(S0,S1, I0[1], I1[1], I2[1], I3[1], R[1]);
mux_4x1 three(S0,S1, I0[2], I1[2], I2[2], I3[2], R[2]);
mux_4x1 four(S0,S1, I0[3], I1[3], I2[3], I3[3], R[3]);
mux_4x1 five(S0,S1, I0[4], I1[4], I2[4], I3[4], R[4]);
mux_4x1 six(S0,S1, I0[5], I1[5], I2[5], I3[5], R[5]);
mux_4x1 seven(S0,S1, I0[6], I1[6], I2[6], I3[6], R[6]);
mux_4x1 eight(S0,S1, I0[7], I1[7], I2[7], I3[7], R[7]);
mux_4x1 nine(S0,S1, I0[8], I1[8], I2[8], I3[8], R[8]);
mux_4x1 ten(S0,S1, I0[9], I1[9], I2[9], I3[9], R[9]);
mux_4x1 eleven(S0,S1, I0[10], I1[10], I2[10], I3[10], R[10]);
mux_4x1 twelve(S0,S1, I0[11], I1[11], I2[11], I3[11], R[11]);
mux_4x1 thirteen(S0,S1, I0[12], I1[12], I2[12], I3[12], R[12]);
mux_4x1 fourteen(S0,S1, I0[13], I1[13], I2[13], I3[13], R[13]);
mux_4x1 fifteen(S0,S1, I0[14], I1[14], I2[14], I3[14], R[14]);
mux_4x1 sixteen(S0,S1, I0[15], I1[15], I2[15], I3[15], R[15]);
mux_4x1 seventeen(S0,S1, I0[16], I1[16], I2[16], I3[16], R[16]);
mux_4x1 eighteen(S0,S1, I0[17], I1[17], I2[17], I3[17], R[17]);
mux_4x1 nineteen(S0,S1, I0[18], I1[18], I2[18], I3[18], R[18]);
mux_4x1 twenty(S0,S1, I0[19], I1[19], I2[19], I3[19], R[19]);
mux_4x1 twentyone(S0,S1, I0[20], I1[20], I2[20], I3[20], R[20]);
mux_4x1 twentytwo(S0,S1, I0[21], I1[21], I2[21], I3[21], R[21]);
mux_4x1 twentythree(S0,S1, I0[22], I1[22], I2[22], I3[22], R[22]);
mux_4x1 twentyfour(S0,S1, I0[23], I1[23], I2[23], I3[23], R[23]);
mux_4x1 twentyfive(S0,S1, I0[24], I1[24], I2[24], I3[24], R[24]);
mux_4x1 twentysix(S0,S1, I0[25], I1[25], I2[25], I3[25], R[25]);
mux_4x1 twentyseven(S0,S1, I0[26], I1[26], I2[26], I3[26], R[26]);
mux_4x1 twentyeight(S0,S1, I0[27], I1[27], I2[27], I3[27], R[27]);
mux_4x1 twentynine(S0,S1, I0[28], I1[28], I2[28], I3[28], R[28]);
mux_4x1 thirty(S0,S1, I0[29], I1[29], I2[29], I3[29], R[29]);
mux_4x1 thirtyone(S0,S1, I0[30], I1[30], I2[30], I3[30], R[30]);
mux_4x1 thirtytwo(S0,S1, I0[31], I1[31], I2[31], I3[31], R[31]);
endmodule